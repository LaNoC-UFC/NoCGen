 
?    Neste trecho será implementado N_ROT arquiteturas, sendo que N_ROT representa o número
?  de roteadores.Cada arquitetura contém uma tabela de roteamento que deve ser utilizado por
?  um roteador.Esta tabela poderá ser baseada em regiões ou não, depende da seleção do usuário.
!
